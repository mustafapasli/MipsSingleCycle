module and_32b(O, A, B);

	input [31:0] A;
	input [31:0] B;

	output [31:0] O;

	and (O[0], A[0], B[0]);
	and (O[1], A[1], B[1]);
	and (O[2], A[2], B[2]);
	and (O[3], A[3], B[3]);
	and (O[4], A[4], B[4]);
	and (O[5], A[5], B[5]);
	and (O[6], A[6], B[6]);
	and (O[7], A[7], B[7]);
	and (O[8], A[8], B[8]);
	and (O[9], A[9], B[9]);
	and (O[10], A[10], B[10]);
	and (O[11], A[11], B[11]);
	and (O[12], A[12], B[12]);
	and (O[13], A[13], B[13]);
	and (O[14], A[14], B[14]);
	and (O[15], A[15], B[15]);
	and (O[16], A[16], B[16]);
	and (O[17], A[17], B[17]);
	and (O[18], A[18], B[18]);
	and (O[19], A[19], B[19]);
	and (O[20], A[20], B[20]);
	and (O[21], A[21], B[21]);
	and (O[22], A[22], B[22]);
	and (O[23], A[23], B[23]);
	and (O[24], A[24], B[24]);
	and (O[25], A[25], B[25]);
	and (O[26], A[26], B[26]);
	and (O[27], A[27], B[27]);
	and (O[28], A[28], B[28]);
	and (O[29], A[29], B[29]);
	and (O[30], A[30], B[30]);
	and (O[31], A[31], B[31]);


endmodule