module nor_32b(O, A, B);

	input [31:0] A;
	input [31:0] B;

	output [31:0] O;

	nor (O[0], A[0], B[0]);
	nor (O[1], A[1], B[1]);
	nor (O[2], A[2], B[2]);
	nor (O[3], A[3], B[3]);
	nor (O[4], A[4], B[4]);
	nor (O[5], A[5], B[5]);
	nor (O[6], A[6], B[6]);
	nor (O[7], A[7], B[7]);
	nor (O[8], A[8], B[8]);
	nor (O[9], A[9], B[9]);
	nor (O[10], A[10], B[10]);
	nor (O[11], A[11], B[11]);
	nor (O[12], A[12], B[12]);
	nor (O[13], A[13], B[13]);
	nor (O[14], A[14], B[14]);
	nor (O[15], A[15], B[15]);
	nor (O[16], A[16], B[16]);
	nor (O[17], A[17], B[17]);
	nor (O[18], A[18], B[18]);
	nor (O[19], A[19], B[19]);
	nor (O[20], A[20], B[20]);
	nor (O[21], A[21], B[21]);
	nor (O[22], A[22], B[22]);
	nor (O[23], A[23], B[23]);
	nor (O[24], A[24], B[24]);
	nor (O[25], A[25], B[25]);
	nor (O[26], A[26], B[26]);
	nor (O[27], A[27], B[27]);
	nor (O[28], A[28], B[28]);
	nor (O[29], A[29], B[29]);
	nor (O[30], A[30], B[30]);
	nor (O[31], A[31], B[31]);


endmodule