`define DELAY 20
module add_32b_testbench();

reg [31:0] A;
reg [31:0] B;
reg C_in;

wire [31:0] O;
wire C_out;

add_32b add32tb (O,C_out, A, B, C_in);

initial begin

C_in = 1'b0;

A = 32'b00000000000000000000000000000011 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000000000000001000100 ; B = 32'b00000000000000000000001000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000100000000000000001 ; B = 32'b00000000100000000000000000000001;
#`DELAY ;
A = 32'b10000000000000000000000000000000 ; B = 32'b10000000000000000000000000000000;
#`DELAY ;
A = 32'b10000010000000000000000000000000 ; B = 32'b10000000000000000000100000000001;
#`DELAY ;
A = 32'b00000000000100000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b10000000010000000000000000000001 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;

C_in = 1'b1;

A = 32'b00000000000000000000000000000011 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000000000000001000100 ; B = 32'b00000000000000000000001000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000100000000000000001 ; B = 32'b00000000100000000000000000000001;
#`DELAY ;
A = 32'b10000000000000000000000000000000 ; B = 32'b10000000000000000000000000000000;
#`DELAY ;
A = 32'b10000010000000000000000000000000 ; B = 32'b10000000000000000000100000000001;
#`DELAY ;
A = 32'b00000000000100000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b10000000010000000000000000000001 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;

end

initial begin

$monitor("time = %2d, A = %10d, B = %10d, R = %10d, C_out = %1b ",$time, A, B, O, C_out);

end

endmodule 