`define DELAY 20
module sub_32b_testbench();

reg [31:0] A;
reg [31:0] B;
reg C_in;

wire [31:0] O;
wire C_out;
wire V;

sub_32b sub32tb (O, V,C_out, A, B, C_in);

initial begin

C_in = 1'b0;

A = 32'b00000000000000000000000000000010 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000010;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000100000000000000001 ; B = 32'b00000000100000000000000000000001;
#`DELAY ;
A = 32'b10000000000000000000000000000001 ; B = 32'b10000000000000000000000000000010;
#`DELAY ;
A = 32'b10000010000000000000000000000000 ; B = 32'b10000000000000000000100000000001;
#`DELAY ;
A = 32'b00000000000100000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b10000000010000000000000000000001 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;

C_in = 1'b1;

A = 32'b00000000000000000000000000000010 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000010;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000100000000000000001 ; B = 32'b00000000100000000000000000000001;
#`DELAY ;
A = 32'b10000000000000000000000000000001 ; B = 32'b10000000000000000000000000000010;
#`DELAY ;
A = 32'b10000010000000000000000000000000 ; B = 32'b10000000000000000000100000000001;
#`DELAY ;
A = 32'b00000000000100000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b10000000010000000000000000000001 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;

end

initial begin

$monitor("time = %2d,C_in = %1b, A = %32b, B = %32b, R = %32b, C_out = %1b, V = %1b ",$time,C_in, A, B, O, C_out, V);

end

endmodule 