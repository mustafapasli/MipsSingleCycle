module or_32b(O, A, B);

	input [31:0] A;
	input [31:0] B;

	output [31:0] O;

	or (O[0], A[0], B[0]);
	or (O[1], A[1], B[1]);
	or (O[2], A[2], B[2]);
	or (O[3], A[3], B[3]);
	or (O[4], A[4], B[4]);
	or (O[5], A[5], B[5]);
	or (O[6], A[6], B[6]);
	or (O[7], A[7], B[7]);
	or (O[8], A[8], B[8]);
	or (O[9], A[9], B[9]);
	or (O[10], A[10], B[10]);
	or (O[11], A[11], B[11]);
	or (O[12], A[12], B[12]);
	or (O[13], A[13], B[13]);
	or (O[14], A[14], B[14]);
	or (O[15], A[15], B[15]);
	or (O[16], A[16], B[16]);
	or (O[17], A[17], B[17]);
	or (O[18], A[18], B[18]);
	or (O[19], A[19], B[19]);
	or (O[20], A[20], B[20]);
	or (O[21], A[21], B[21]);
	or (O[22], A[22], B[22]);
	or (O[23], A[23], B[23]);
	or (O[24], A[24], B[24]);
	or (O[25], A[25], B[25]);
	or (O[26], A[26], B[26]);
	or (O[27], A[27], B[27]);
	or (O[28], A[28], B[28]);
	or (O[29], A[29], B[29]);
	or (O[30], A[30], B[30]);
	or (O[31], A[31], B[31]);


endmodule