`define DELAY 20
module and_32b_testbench();

reg [31:0] A;
reg [31:0] B;

wire [31:0] R;

and_32b and32tb (R, A, B);

initial begin

A = 32'b00000000000000000000000000000000 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000000000000000000000 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000000 ; B = 32'b10000000000000000000000000000000;
#`DELAY ;
A = 32'b10000000000000000000000000000000 ; B = 32'b10000000000000000000000000000001;
#`DELAY ;
A = 32'b00000000000000000000000000000001 ; B = 32'b00000000000000000000000000000000;
#`DELAY ;
A = 32'b10000000000000000000000000000001 ; B = 32'b00000000000000000000000000000001;
#`DELAY ;

end

initial begin

$monitor("time = %2d, A = %32b, B = %32b, R = %32b",$time, A, B, R);

end

endmodule 