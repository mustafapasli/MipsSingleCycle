`define DELAY 20
module shift_32b_testbench();

reg D; 

reg [31:0] A,  B;

wire [31:0] O;

shift_32b s32btb (O, A, B, D); //  D> direction, F> false=0

initial begin

A = 32'b10000000000000100000000000000001;

B = 32'b00000000000000000000000000000001; D = 1'b0;
#`DELAY;
B = 32'b00000000000000000000000000000001; D = 1'b1;
#`DELAY;
B = 32'b00000000000000000000000000000011; D = 1'b0;
#`DELAY;
B = 32'b00000000000000000000000000000011; D = 1'b1; 
#`DELAY;
B = 32'b00000000000000000000000000000111; D = 1'b0;
#`DELAY;
B = 32'b00000000000000000000000000000111; D = 1'b1;
#`DELAY;
B = 32'b00000000000000000000000000001111; D = 1'b0;
#`DELAY;
B = 32'b00000000000000000000000000001111; D = 1'b1; 
#`DELAY;
B = 32'b00000000000010000000000000000000; D = 1'b0;
#`DELAY;
B = 32'b00000000000010000000000000000000; D = 1'b1; 
#`DELAY;


end

initial begin

$monitor("time = %2d, A = %32b, B = %32b, D = %1b, O = %32b ",$time,A, B, D, O);

end

endmodule